module keyboard(S);